----------------------------------------------------------------------------------
-- Company: Univesidad de Zaragoza
-- Engineer: Javier Resano/Jose Luis Briz
-- 
-- Create Date:    10:38:16 27/12/2024 
-- Design Name: 
-- Module Name:    memoriaRAM_I - Behavioral 

-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_unsigned.all;
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity memoriaRAM_I is port (
		  	CLK : in std_logic;
		  	ADDR : in std_logic_vector (31 downto 0); --Dir 
        	Din : in std_logic_vector (31 downto 0);--entrada de datos para el puerto de escritura
        	WE : in std_logic;		-- write enable	
		  	RE : in std_logic;		-- read enable		  
		  	Dout : out std_logic_vector (31 downto 0));
end memoriaRAM_I;

--************************************************************************************************************
-- Instruction memory file loaded with various tests.
-- IMPORTANT: There can only be one uncommented test. 
-- To run a test, uncomment it, and comment on the rest.
--************************************************************************************************************

architecture Behavioral of memoriaRAM_I is
type RamType is array(0 to 127) of std_logic_vector(31 downto 0);
--------------------------------------------------------------------------------------------------------------------------------
-- Instruction Memory Map
-- From Word 0 to 3: Exception Vector Table: (@ of the exception routines)
-- 		@0: reset
-- 		@4: IRQ
-- 		@8: Data Abort
-- 		@C: UNDEF
-- From Word 4  (@010): .CODE (code of the application to execute)
-- From Word 64 (@100): RTI (code for the IRQ)
-- From Word 96 (@180): Data abort (code for the Data Abort exception)
-- From Word 112(@1C0): UNDEF (code for the UNDEF exception)
--------------------------------------------------------------------------------------------------------------------------------


--------------------------------------------------------------------------------------------------------------------------------
-- TESTBENCH 1: Delayed SYSTEM 
-- Delayed_code including nops to eliminate data and control hazards. 
-- It loops infinitely in case of IRQ, undef, or abort exceptions.
-- Code overview: MEM[0]= MEM[0] + MEM[4]; while(1);//MEM[0]=256+1
-- Reset: beq R1, R1, INI; 
-- Ini: LW  R31, 0(R0); 
-- Main: LW  R1, 0(R0); LW  R2, 4(R0); NOP; NOP; ADD R3, R1, R2; NOP; NOP; SW  R3, 0(R0); end: beq r0, r0, end; NOP
-- It should work on the initial processor. 
-- NEXT STEPS: 
-- 1) After designing the hazard-detection and fordwarding units, remove the unnecessary nops and check that it still works.
-- 2) Replace the 4 instructions in the loop with a lw_inc and check that you get the same result. 
--------------------------------------------------------------------------------------------------------------------------------
--signal RAM : RamType := (  			X"10210003", X"00000000", X"00000000", X"00000000", X"081F0000", X"08010000", X"08020004", X"00000000", --word 0,1,...
--									X"00000000", X"04221800", X"00000000", X"00000000", X"0C030008", X"1000FFFF", X"00000000", X"00000000", --word 8,9,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 16,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 24,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 32,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 40,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 48,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 56,...
--									X"1000FFFF", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 64,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",--word 72,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 80,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 88,...
--									X"1000FFFF", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 96,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 104,...
--									X"1000FFFF", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 112,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000");--word 120,...										
--														
--------------------------------------------------------------------------------------------------------------------------------
-- TESTBENCH 2: for IRQ and mutual exclusion between IRQ and main with LW_inc
-- Described in detail in Testbench_IRQ_2025
--------------------------------------------------------------------------------------------------------------------------------
-- signal RAM : RamType := ( X"10210003", X"1021003E", X"1021005D", X"1021006C", X"081F0000", X"40010020", X"08020024", X"10220001",--word 0,1,...
-- 									X"1021FFFD", X"08010008", X"0C017004", X"0C027004", X"40010024", X"1021FFF7", X"00000000", X"00000000", --word 8,9,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 16,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 24,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 32,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 40,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 48,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 56,...
--									X"0FE10000", X"0FE20004", X"08C10008", X"07E1F800", X"08010028", X"08020024", X"10220001", X"10210006", --word 64,...
--									X"08010000", X"0C017004", X"0C027004", X"40010020", X"0C010028", X"40010024", X"08010004", X"0CC17008", --word 72,...
--									X"08010008", X"07E1F801", X"0BE10000", X"0BE20004", X"20000000", X"08C17FFF", X"00000000", X"00000000",--word 80,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 88,...
--									X"08C10014", X"0CC67004", X"0CC17004", X"20000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 96,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 104,...
--									X"08C1001C", X"0CC17004", X"1000FFFF", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 112,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000");--word 120,...
									
								
--------------------------------------------------------------------------------------------------------------------------------
-- TESTBENCH 3: DATA ABORT 1
-- Unaligned memory access: 08010003 = LW R1, 3(R0)
-- Produces an abort and we jump to word 96 which outputs the code 0x00000AB0 and enters an infinite loop: 1000FFFF = BEQ r0,r0,-1
-- There is an RTE after the loop which, if everything is well managed, will never be executed.
--------------------------------------------------------------------------------------------------------------------------------
 --signal RAM : RamType := (  			X"10210003", X"1021003E", X"1021005D", X"1021006C", X"08010003", X"00000000", X"00000000", X"00000000", --word 0,1,...
-- 									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 8,9,...
-- 									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 16,...
-- 									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 24,...
-- 									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 32,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 40,...
 --									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 48,...
 --									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 56,...
 --									X"0FE10000", X"0FE20004", X"08C10008", X"07E1F800", X"08C2000C", X"08C10004", X"04221000", X"0CC27004", --word 64,...
 --									X"0CC2000C", X"0CC17008", X"08C10008", X"07E1F801", X"0BE10000", X"0BE20004", X"20000000", X"08C17FFF",--word 72,...
 --									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 80,...
 --									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 88,...
 --									X"08C10014", X"0CC17004", X"1000FFFF", X"20000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 96,...
 --									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 104,...
 --									X"08C1001C", X"0CC17004", X"1000FFFF", X"20000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 112,...
 --									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000");--word 120,...
 --									
--------------------------------------------------------------------------------------------------------------------------------
-- TESTBENCH 4: DATA ABORT 2
-- Access to out-of-range address: 08017ffC = LW R1, 32767(R0)
-- Produces an abort and we jump to word 96 which outputs the code 0x00000AB0 and enters an infinite loop: 1000FFFF = BEQ r0,r0,-1
-- There is an RTE after the loop which, if everything is well managed, will never be executed.
--------------------------------------------------------------------------------------------------------------------------------
-- signal RAM : RamType := (  		X"10210003", X"1021003E", X"1021005D", X"1021006C", X"08017ffC", X"00000000", X"00000000", X"00000000", --word 0,1,...
-- 									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 8,9,...
-- 									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 16,...
-- 									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 24,...
-- 									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 32,...
-- 									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 40,...
-- 									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 48,...
-- 									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 56,...
-- 									X"0FE10000", X"0FE20004", X"08C10008", X"07E1F800", X"08C2000C", X"08C10004", X"04221000", X"0CC27004", --word 64,...
-- 									X"0CC2000C", X"0CC17008", X"08C10008", X"07E1F801", X"0BE10000", X"0BE20004", X"20000000", X"08C17FFF",--word 72,...
-- 									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 80,...
-- 									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 88,...
-- 									X"08C10014", X"0CC17004", X"1000FFFF", X"20000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 96,...
-- 									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 104,...
-- 									X"08C1001C", X"0CC17004", X"1000FFFF", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 112,...
-- 									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000");--word 120,...
-- 									
--------------------------------------------------------------------------------------------------------------------------------
-- TESTBENCH 5: UNDEF
-- Instruction with incorrect code: FFFFFFFF = �?
-- Produces an UNDEF and the execution jumps to word 112 which outputs the code 0x0BAD0C0D and enters an infinite loop: 1000FFFF = BEQ r0,r0,-1
-- There is an RTE after the loop which, if everything is well managed, will never be executed.
--------------------------------------------------------------------------------------------------------------------------------
-- signal RAM : RamType := (  		X"10210003", X"1021003E", X"1021005D", X"1021006C", X"FFFFFFFF", X"00000000", X"00000000", X"00000000", --word 0,1,...
-- 									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 8,9,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 16,...
-- 									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 24,....
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 32,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 40,...
-- 									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 48,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 56,...
--									X"0FE10000", X"0FE20004", X"08C10008", X"07E1F800", X"08C2000C", X"08C10004", X"04221000", X"0CC27004", --word 64,...
--									X"0CC2000C", X"0CC17008", X"08C10008", X"07E1F801", X"0BE10000", X"0BE20004", X"20000000", X"08C17FFF",--word 72,...
-- 									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 80,...
-- 									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 88,...
-- 									X"08C10014", X"0CC17004", X"1000FFFF", X"20000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 96,...
-- 									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 104,...
-- 									X"08C1001C", X"0CC17004", X"1000FFFF", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 112,...
-- 									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000");--word 120,...

-----------------------------------------------------------------------------------------------------------------------------

--------------------------------------------------------------------------------------------------------------------------------
-- TESTBENCH 6: Prueba pr3
-- Probamos si funciona el programa de la p?actica 3, es decir probamos el funcionamiento de las instrucciones
-- JAL y RET, al igual que un caso de forwarding.
--------------------------------------------------------------------------------------------------------------------------------
-- signal RAM : RamType := (  		X"10000003", X"10000007", X"10000006", X"10000005", X"08010018", X"0802001C", X"08030020", X"14070002", X"0C050014", X"1000FFFF", X"10230004", X"08260000", --word 0,1,...
--									X"04220800", X"04A62800", X"1000FFFB", X"18E70000",  --word 8,9,...
--									X"08010004", X"0CC17008", X"20000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 16,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 24,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 32,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 40,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 48,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 56,...
--									X"0FE10000", X"0FE20004", X"08C10008", X"07E1F800", X"08C2000C", X"08C10004", X"04221000", X"0CC27004", --word 64,...
--									X"0CC2000C", X"0CC17008", X"08C10008", X"07E1F801", X"0BE10000", X"0BE20004", X"20000000", X"08C17FFF",--word 72,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 80,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 88,...
--									X"08C10014", X"0CC17004", X"1000FFFF", X"20000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 96,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 104,...
--									X"08C1001C", X"0CC17004", X"1000FFFF", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 112,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000");--word 120,...
-----------------------------------------------------------------------------------------------------------------------------

--------------------------------------------------------------------------------------------------------------------------------
-- TESTBENCH 7: Prueba adelantamiento operandos distancia 1-2 y paradas si son necesarias.
-- Probamos funcionan las paradas a distancia 1 con mismos operados, adelantamiento a de operandos a distancias
-- 1 y 2 de las operaciones.
--------------------------------------------------------------------------------------------------------------------------------
-- signal RAM : RamType := (  		X"40010014", X"40010014", X"04210800", X"0C01001C", X"04411000", X"04221800", X"0C030018", X"10230005", --word 0,1,...
-- 								X"04231801", X"04431800", X"10000002", X"00000000", X"00000000", X"1000FFFF", X"10000006", X"10000005",  --word 8,9,...
-- 								X"08010004", X"0CC17008", X"08040020", X"18800000", X"08040024", X"00000000", X"18A00000", X"20000000", --word 16,...
-- 								X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 24,...
-- 								X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 32,...
-- 								X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 40,...
-- 								X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 48,...
-- 								X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 56,...
-- 								X"0FE10000", X"0FE20004", X"08C10008", X"07E1F800", X"08C2000C", X"08C10004", X"04221000", X"0CC27004", --word 64,...
-- 								X"0CC2000C", X"0CC17008", X"08C10008", X"07E1F801", X"0BE10000", X"0BE20004", X"20000000", X"08C17FFF",--word 72,...
-- 								X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 80,...
-- 								X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 88,...
-- 								X"08C10014", X"0CC17004", X"1000FFFF", X"20000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 96,...
-- 								X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 104,...
-- 								X"08C1001C", X"0CC17004", X"1000FFFF", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 112,...
-- 								X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000");--word 120,...
-----------------------------------------------------------------------------------------------------------------------------

--------------------------------------------------------------------------------------------------------------------------------
-- TESTBENCH 1 P2: Unit test (1)
--------------------------------------------------------------------------------------------------------------------------------
---signal RAM : RamType := (
--    X"08010060", X"0C020060", X"0C0200A0", X"080300A0", X"08040070", X"08050074", X"08060078", X"00000000", --word 0,1,...
--    X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 8,9,...
--   X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 16,...
 --   X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 24,...
 --   X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 32,...
   -- X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 40,...
--    X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 48,...
--    X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 56,...
--    X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 64,...
--    X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 72,...
--    X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 80,...
--    X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 88,...
--    X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 96,...
--    X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 104,...
--    X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 112,...
--    X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000");--word 120,...

--------------------------------------------------------------------------------------------------------------------------------
-- TESTBENCH ERROR P2: Unit test (1)
--------------------------------------------------------------------------------------------------------------------------------  
-- signal RAM : RamType := (
--     X"10210003", X"1021000F", X"10210011", X"10210016", X"08020004", X"08030008", X"0C430004", X"0803000C", --word 0,1,...
--     X"0C430008", X"40040041", X"08650000", X"0C05000C", X"08060200", X"080601FC", X"0C060020", X"0C660000", --word 8,9,...
--     X"1000FFFF", X"08010000", X"0C017008", X"20000000", X"08410004", X"0C017004", X"08410008", X"08210000", --word 16,...
--     X"0C010030", X"20000000", X"08010010", X"0C017004", X"1000FFFC", X"00000000", X"00000000", X"00000000", --word 24,...
--     X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 32,...
--     X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 40,...
--     X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 48,...
--     X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 56,...
--     X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 64,...
--     X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 72,...
--     X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 80,...
--     X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 88,...
--     X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 96,...
--     X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 104,...
--     X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 112,...
--     X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000");--word 120,...
--------------------------------------------------------------------------------------------------------------------------------
-- TESTBENCH P2: Huge Unit Test 1
--------------------------------------------------------------------------------------------------------------------------------
-- signal RAM : RamType := (
--  X"04000000", X"08010060", X"08010064", X"08020020", X"08020028", X"0C010010", X"08030014", X"0C030010", --word 0,1,...
--  X"0C020050", X"08020050", X"08040054", X"0801006C", X"08020024", X"080500A0", X"40080060", X"080600E0", --word 8,9,...
--  X"400600E0", X"400500A4", X"40040040", X"080600E4", X"0C060090", X"0C0700D0", X"0C0100A0", X"0C0100E0", --word 16,...
--  X"0C020094", X"0C0200D8", X"08010090", X"08010094", X"08010098", X"0801009C", X"08010000", X"08020040", --word 24,...
--  X"40010080", X"08010000", X"08010080", X"08010000", X"0C010044", X"0C010090", X"00000000", X"00000000", --word 32,...
--  X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 40,...
--  X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 48,...
--  X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 56,...
--  X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 64,...
--  X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 72,...
--  X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 80,...
--  X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 88,...
--  X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 96,...
--  X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 104,...
--  X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 112,...
--  X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000");--word 120,...
--------------------------------------------------------------------------------------------------------------------------------
-- TESTBENCH P2: Huge Unit Test 2
--------------------------------------------------------------------------------------------------------------------------------
--signal RAM : RamType := (
--    X"08000000", X"0801000C", X"0C010010", X"08010010", X"40010014", X"0BE20004", X"0FE10004", X"0FE10010", --word 0,1,...
--    X"0FE10050", X"0BE30090", X"0BE400D0", X"0FE10090", X"0FE30090", X"0FE40090", X"43E50010", X"0BE30090", --word 8,9,...
--    X"0FE47000", X"0BE47000", X"0FE37004", X"0BE47004", X"0FE27008", X"0BE47008", X"00000000", X"00000000", --word 16,...
--    X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 24,...
--    X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 32,...
--    X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 40,...
--    X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 48,...
--    X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 56,...
--    X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 64,...
--    X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 72,...
--    X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 80,...
--    X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 88,...
--    X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 96,...
--    X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 104,...
--    X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 112,...
--    X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000");--word 120,...
-----------------------------------------------------------------------
-- PARA ANÁLISIS DE LATENCIAS
----------------------------------------------------------------------------
-- signal RAM : RamType := (
--     X"0C010000", X"40010000", X"40010000", X"0C010000", X"08020004", X"08430004", X"04611800", X"0C430004", --word 0,1,...
--     X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 8,9,...
--     X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 16,...
--     X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 24,...
--     X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 32,...
--     X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 40,...
--     X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 48,...
--     X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 56,...
--     X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 64,...
--     X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 72,...
--     X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 80,...
--     X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 88,...
--     X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 96,...
--     X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 104,...
--     X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 112,...
--     X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000");--word 120,...
-----------------------------------------------------------------------
-- RAM PARA ETHICAL HACKING
----------------------------------------------------------------------------
-- signal RAM : RamType := (
--     X"08000000", X"08010004", X"08020008", X"0803000C", X"04632000", X"04842000", X"04052800", X"04263000", --word 0,1,...
--     X"04473800", X"04684000", X"0D200000", X"0D200040", X"0D200080", X"0D2000C0", X"0D210010", X"0D210050", --word 8,9,...
--     X"0D210090", X"0D2100D0", X"0D220020", X"0D220060", X"0D2200A0", X"0D2200E0", X"0D230030", X"0D230070", --word 16,...
--     X"0D2300B0", X"0D2300F0", X"04050000", X"04260800", X"04471000", X"04681800", X"04852001", X"11240001", --word 24,...
--     X"1000FFE9", X"09200000", X"09210040", X"09220080", X"092300C0", X"04010000", X"04020000", X"04030000", --word 32,...
--     X"0D200000", X"09200010", X"09210050", X"09220090", X"092300D0", X"04010000", X"04020000", X"04030000", --word 40,...
--     X"0D200040", X"09200020", X"09210060", X"092200A0", X"092300E0", X"04010000", X"04020000", X"04030000", --word 48,...
--     X"0D200080", X"09200030", X"09210070", X"092200B0", X"092300F0", X"04010000", X"04020000", X"04030000", --word 56,...
--     X"0D2000C0", X"1000FFFF", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 64,...
--     X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 72,...
--     X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 80,...
--     X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 88,...
--     X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 96,...
--     X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 104,...
--     X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 112,...
--     X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000");--word 120,...
-----------------------------------------------------------------------
-- RAM PARA TEST INTEGRADO
-----------------------------------------------------------------------
signal RAM : RamType := (
    X"04000000", X"04007000", X"04007800", X"080A00FC", X"080B010C", X"080C0108", X"056B6800", X"05AD6800", --word 0,1,...
    X"04000800", X"08020100", X"08030104", X"08240000", X"08450000", X"04853000", X"08240004", X"08450004", --word 8,9,...
    X"04853800", X"08240004", X"08450004", X"04854000", X"08240004", X"08450004", X"04854800", X"0C660000", --word 16,...
    X"0C670004", X"0C680008", X"0C69000C", X"042C0800", X"044C1000", X"046C1800", X"05EB7800", X"11AF0001", --word 24,...
    X"1000FFEA", X"04007800", X"08010104", X"08030110", X"08240000", X"04842800", X"08240004", X"04843000", --word 32,...
    X"08240008", X"04843800", X"0824000C", X"04844000", X"0C250000", X"0C260004", X"0C270008", X"0C28000C", --word 40,...
    X"042C0800", X"05EB7800", X"11AF0001", X"1000FFF0", X"08020100", X"40440000", X"40440010", X"40440020", --word 48,...
    X"40440030", X"04007800", X"04000800", X"08020100", X"08030114", X"08240000", X"08450000", X"04853000", --word 56,...
    X"08240004", X"08450004", X"04853800", X"08240004", X"08450004", X"04854000", X"08240004", X"08450004", --word 64,...
    X"04854800", X"0C660000", X"0C670004", X"0C680008", X"0C69000C", X"042C0800", X"044C1000", X"046C1800", --word 72,...
    X"05EB7800", X"11AF0001", X"1000FFEA", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 80,...
    X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 88,...
    X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 96,...
    X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 104,...
    X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 112,...
    X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000");--word 120,...
signal dir_7:  std_logic_vector(6 downto 0); 
begin
 
 dir_7 <= ADDR(8 downto 2); -- As the memory is 128 words we do not use the full address but only 7 bits. As bytes are addressed, but we give words we do not use the 2 least significant bits.
 process (CLK)
    begin
        if (CLK'event and CLK = '1') then
            if (WE = '1') then -- It is written only if WE is 1
                RAM(conv_integer(dir_7)) <= Din;
            end if;
        end if;
    end process;

    Dout <= RAM(conv_integer(dir_7)) when (RE='1') else "00000000000000000000000000000000"; -- It is only read if RE is 1

end Behavioral;


